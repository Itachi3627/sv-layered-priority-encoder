class driver;
    virtual intf.driver vif;
    mailbox #(transaction) gen2drv;
    transaction trans;

    function new(virtual intf.driver vif, mailbox #(transaction) g2d);
        this.vif = vif;
        this.gen2drv = g2d;
    endfunction

  task run();
        $display("[DRIVER] Starting driver");  
        forever begin 
            gen2drv.get(trans);
            driver_trans(trans);
        end
    endtask

    task driver_trans(transaction trans);
        vif.req =  trans.req;
        #5;
        ->vif.sample_enable;
        #5;
    endtask

endclass